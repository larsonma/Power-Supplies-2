****************************************************
* Filename: lab4.cir
* Author: 	larsonma@msoe.edu <Mitchell Larson>
* Date:		March 27th 2018
* Provides:
*	- DC power supply design simulation
*	- VS = 120 VRMS - main voltage
*	- V2 = 12 VRMS - voltage after transformer
*	- Vr = 0.5V	
*	- RL = 1000 Ohm
*	- Vo = 5 VDC
*	- VM = 12 VRMS = 16.973V - 1.4V
****************************************************

*** Semiconductor Model ***
* - Modeled after the DB101 Full Bridge Rectifier
.model DB101 D(Is=7.3155p, Bv = 50, N=1.5, Rs=0.05)


*** US Power Thevenin ***
VS 1 0 SIN(0,170,60)
RP 1 2 0.1

*** Transformer modeled as inductors ***
L1 2 0 10m
L2 3 5 100u
K1 L1 L2 0.99

*** Joining isolated circuits to common ground for PSPICE simulation ***
RSIM 5 0 1000MEG

*** Full-wave bridge rectifier ***
D1 3 4 DB101
D2 0 5 DB101
D3 5 4 DB101
D4 0 3 DB101

*** Filter capacitance ***
C1 4 0 2.60m

*** Load resistance ***
RL 4 0 1000

*** Control Statements ***
.tran 0.001m 33.34m

*** request oscope ***
.probe

.end